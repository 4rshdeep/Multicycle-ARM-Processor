entity data_path is
  port (
	clock
  ) ;
end entity ; 